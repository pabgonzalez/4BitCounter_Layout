magic
tech sky130A
magscale 1 2
timestamp 1710021771
<< nwell >>
rect -36 -794 2763 649
<< poly >>
rect -94 -709 -61 1767
rect 1771 -830 1994 -800
rect 2098 -825 2226 -811
rect -10 -922 114 -892
rect -10 -1339 25 -922
rect 1857 -1269 1887 -830
rect 2073 -841 2226 -825
rect 2196 -1329 2226 -841
rect 2758 -1229 2793 2100
rect 2757 -1336 2793 -1229
<< metal1 >>
rect 2427 2071 2757 2106
rect -90 1738 951 1771
rect -90 1737 10 1738
rect -75 -680 -6 -675
rect -75 -713 75 -680
rect -75 -714 -6 -713
rect 2112 -718 2369 -716
rect 2026 -750 2369 -718
rect 2026 -752 2282 -750
rect -9 -1307 2228 -1305
rect -9 -1339 2793 -1307
rect 2193 -1341 2793 -1339
use dffc  dffc_0 ../dffc
timestamp 1710021771
transform 1 0 900 0 1 1174
box -900 -1174 1816 1067
use inverter  inverter_1 ../inverter
timestamp 1710021771
transform 1 0 1731 0 1 -1783
box 474 522 794 1585
use nand  nand_1 ../nand
timestamp 1710021771
transform 1 0 1889 0 1 -1261
box 0 0 320 1063
use via_m1_p#1  via_m1_p_0 ../via_m1_p
timestamp 1646951168
transform 1 0 -27 0 1 -1357
box 0 0 68 68
use via_m1_p#1  via_m1_p_1
timestamp 1646951168
transform 1 0 2742 0 1 -1357
box 0 0 68 68
use via_m1_p#1  via_m1_p_2
timestamp 1646951168
transform 1 0 2177 0 1 -1357
box 0 0 68 68
use via_m1_p#1  via_m1_p_3
timestamp 1646951168
transform 1 0 -112 0 1 1716
box 0 0 68 68
use via_m1_p#1  via_m1_p_4
timestamp 1646951168
transform 1 0 -113 0 1 -726
box 0 0 68 68
use via_m1_p#1  via_m1_p_5
timestamp 1646951168
transform 1 0 2332 0 1 -768
box 0 0 68 68
use via_m1_p#1  via_m1_p_13
timestamp 1646951168
transform -1 0 2811 0 -1 2117
box 0 0 68 68
use xor  xor_1 ../xor
timestamp 1710021771
transform -1 0 1559 0 1 -1272
box -323 13 1551 1078
<< labels >>
rlabel poly 1857 -1269 1887 -800 1 ce
rlabel space 2664 2 2700 1650 1 clr
rlabel space 252 1374 282 1994 1 clk
rlabel space 2758 -1336 2793 2117 1 Q
rlabel space 2474 -1056 2510 -462 1 sout
<< end >>
