magic
tech sky130A
magscale 1 2
timestamp 1709941173
<< poly >>
rect 622 728 652 1320
rect 744 746 778 1304
<< metal1 >>
rect 494 1504 776 1560
rect 576 1424 610 1504
rect 664 1304 698 1346
rect 664 1270 746 1304
rect 664 746 746 780
rect 664 692 698 746
rect 576 578 610 654
rect 494 522 776 578
use grid  grid_0 ../grid
timestamp 1678218586
transform 1 0 535 0 1 532
box -61 -10 259 1053
use sky130_fd_pr__nfet_01v8_SKHSUU  sky130_fd_pr__nfet_01v8_SKHSUU_0
timestamp 1709668861
transform 1 0 637 0 1 673
box -73 -71 73 71
use sky130_fd_pr__pfet_01v8_52DS5B  sky130_fd_pr__pfet_01v8_52DS5B_0
timestamp 1709668672
transform 1 0 637 0 1 1383
box -109 -107 109 107
use via_m1_p  via_m1_p_0 ../via_m1_p
timestamp 1646951168
transform 1 0 726 0 1 728
box 0 0 68 68
use via_m1_p  via_m1_p_2
timestamp 1646951168
transform 1 0 726 0 1 1252
box 0 0 68 68
<< labels >>
rlabel poly 622 728 652 1320 1 in
rlabel metal1 494 1504 776 1560 1 vdd
rlabel metal1 494 522 776 578 1 vss
rlabel space 744 728 778 1320 1 out
<< end >>
