magic
tech sky130A
magscale 1 2
timestamp 1709822015
<< poly >>
rect 188 942 478 976
rect 446 432 478 942
rect 102 196 132 304
rect 534 196 564 246
rect 102 162 564 196
<< metal1 >>
rect 56 914 90 986
rect 300 476 522 504
rect 232 282 266 334
rect 300 282 334 476
rect 488 406 522 476
rect 232 252 334 282
rect 400 54 434 272
rect 576 40 610 268
use grid  grid_0 grid
timestamp 1678218586
transform 1 0 381 0 1 10
box -61 -10 259 1053
use grid  grid_1
timestamp 1678218586
transform 1 0 61 0 1 10
box -61 -10 259 1053
use sky130_fd_pr__nfet_01v8_NDWVGB  sky130_fd_pr__nfet_01v8_NDWVGB_1
timestamp 1709815372
transform 1 0 461 0 1 340
box -73 -101 73 101
use sky130_fd_pr__nfet_01v8_NDWVGB  sky130_fd_pr__nfet_01v8_NDWVGB_2
timestamp 1709815372
transform 1 0 549 0 1 340
box -73 -101 73 101
use sky130_fd_pr__pfet_01v8_5EUKDE  sky130_fd_pr__pfet_01v8_5EUKDE_0
timestamp 1709817887
transform 1 0 205 0 1 625
box -109 -362 109 362
use sky130_fd_pr__pfet_01v8_5EUKDE  sky130_fd_pr__pfet_01v8_5EUKDE_1
timestamp 1709817887
transform 1 0 117 0 1 625
box -109 -362 109 362
<< labels >>
rlabel metal1 232 252 334 282 1 Z
rlabel poly 102 162 564 196 1 B
rlabel poly 446 432 478 976 1 A
<< end >>
