** sch_path: /foss/designs/tests/test1_4BitCounter.sch
**.subckt test1_4BitCounter
x2 avdd1p8 net1 q0 avss1p8 inverter
V4 avss1p8 GND DC{vss}
V5 avdd1p8 avss1p8 DC{vdd}
V6 ce avss1p8 PULSE(0 {vdd} {Tclk/4} 1p 1p {22*Tclk} {25*Tclk}) DC 0 AC 0
C1 net1 avss1p8 1p m=1
V1 clk avss1p8 PULSE({vdd} 0 0.0 1p 1p {Tclk/2} {Tclk}) DC 0 AC 0
V2 clr avss1p8 PULSE(0 {vdd} {-Tclk/2} 1p 1p {Tclk*2} {Tclk*30}) DC 0 AC 0
x1 q2 q1 q0 q3 clr clk ce avdd1p8 avss1p8 4BitCounter
x3 avdd1p8 net2 q1 avss1p8 inverter
C2 net2 avss1p8 1p m=1
x4 avdd1p8 net3 q2 avss1p8 inverter
C3 net3 avss1p8 1p m=1
x5 avdd1p8 net4 q3 avss1p8 inverter
C4 net4 avss1p8 1p m=1
**** begin user architecture code


* Circuit Parameters
.param vdd = 1.8
.param vss = 0.0
.param Tclk = 15n
.options TEMP = 65.0

* Include Models
.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice TT

* OP Parameters & Singals to save
.save all

* Simulations
.control
  tran 0.01u 1u
  setplot tran1
  plot clr ce+2 v(q0)+4 v(q1)+6 v(q2)+8 v(q3)+10 clk+12
reset
.endc

.end


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/inverter.sym # of pins=4
** sym_path: /foss/designs/inverter.sym
** sch_path: /foss/designs/inverter.sch
.subckt inverter vdd out in vss
*.iopin out
*.iopin vss
*.iopin vdd
*.iopin in
XM2 out in vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 out in vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=0.45 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /foss/designs/4BitCounter.sym # of pins=9
** sym_path: /foss/designs/4BitCounter.sym
** sch_path: /foss/designs/4BitCounter.sch
.subckt 4BitCounter q2 q1 q0 q3 clr clk ce vdd vss
*.iopin ce
*.iopin clk
*.iopin clr
*.iopin q0
*.iopin q1
*.iopin q2
*.iopin q3
*.iopin vss
*.iopin vdd
x1 clr q0 clk ce vdd vss net1 1BitCounter
x2 clr q1 clk net1 vdd vss net2 1BitCounter
x3 clr q2 clk net2 vdd vss net3 1BitCounter
x4 clr q3 clk net3 vdd vss net4 1BitCounter
.ends


* expanding   symbol:  /foss/designs/1BitCounter.sym # of pins=7
** sym_path: /foss/designs/1BitCounter.sym
** sch_path: /foss/designs/1BitCounter.sch
.subckt 1BitCounter clr Q clk ce vdd vss sout
*.iopin clk
*.iopin sout
*.iopin ce
*.iopin clr
*.iopin vdd
*.iopin vss
*.iopin Q
x1 vdd ce sout Q vss and
x2 vdd net1 ce Q vss xor
x3 Q net1 clk clr vss vdd dffc
.ends


* expanding   symbol:  /foss/designs/and.sym # of pins=5
** sym_path: /foss/designs/and.sym
** sch_path: /foss/designs/and.sch
.subckt and vdd A Z B vss
*.iopin Z
*.iopin A
*.iopin B
*.iopin vdd
*.iopin vss
x1 vdd net1 A B vss nand
x2 vdd Z net1 vss inverter
.ends


* expanding   symbol:  /foss/designs/xor.sym # of pins=5
** sym_path: /foss/designs/xor.sym
** sch_path: /foss/designs/xor.sch
.subckt xor vdd Z A B vss
*.iopin A
*.iopin B
*.iopin vdd
*.iopin Z
*.iopin vss
XM6 net1 Bb vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 Z Ab net1 vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 Z A net2 vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 net2 B vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM0 net3 Bb vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 net4 Ab vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Z A net3 vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 Z B net4 vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
x1 vdd Ab A vss inverter
x2 vdd Bb B vss inverter
.ends


* expanding   symbol:  /foss/designs/dffc.sym # of pins=6
** sym_path: /foss/designs/dffc.sym
** sch_path: /foss/designs/dffc.sch
.subckt dffc Q D clk clr vss vdd
*.iopin clk
*.iopin clr
*.iopin vss
*.iopin vdd
*.iopin D
*.iopin Q
x1 vdd n_clk clk vss inverter
x2 vdd net4 net1 vss inverter
x3 vdd Qb Q vss inverter
x4 D p_clk n_clk net1 vss vdd tg
x8 vdd Q clr net3 vss nor
x9 vdd net2 clr net4 vss nor
x5 net2 n_clk p_clk net1 vss vdd tg
x6 net4 n_clk p_clk net3 vss vdd tg
x7 Qb p_clk n_clk net3 vss vdd tg
x10 vdd p_clk n_clk vss inverter
.ends


* expanding   symbol:  /foss/designs/nand.sym # of pins=5
** sym_path: /foss/designs/nand.sym
** sch_path: /foss/designs/nand.sch
.subckt nand vdd Z A B vss
*.iopin B
*.iopin A
*.iopin vdd
*.iopin Z
*.iopin vss
XM1 net1 B vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Z A net1 vss sky130_fd_pr__nfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 Z A vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 Z B vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /foss/designs/tg.sym # of pins=6
** sym_path: /foss/designs/tg.sym
** sch_path: /foss/designs/tg.sch
.subckt tg vin enb en vout vss vdd
*.iopin vin
*.iopin vout
*.iopin enb
*.iopin en
*.iopin vss
*.iopin vdd
XM1 vin en vout vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.75 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 vout enb vin vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /foss/designs/nor.sym # of pins=5
** sym_path: /foss/designs/nor.sym
** sch_path: /foss/designs/nor.sch
.subckt nor vdd Z A B vss
*.iopin A
*.iopin B
*.iopin vdd
*.iopin Z
*.iopin vss
XM1 Z A vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.75 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 B vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 Z B vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=0.75 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 Z A net1 vdd sky130_fd_pr__pfet_01v8 L=0.15 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
