** sch_path: /foss/designs/sch/tests/test1_4BitCounter.sch
**.subckt test1_4BitCounter
*  x2 -  inverter  IS MISSING !!!!
V4 avss1p8 GND DC{vss}
V5 avdd1p8 avss1p8 DC{vdd}
V6 ce avss1p8 PULSE(0 {vdd} {Tclk/4} 1p 1p {22*Tclk} {25*Tclk}) DC 0 AC 0
C1 net1 avss1p8 1p m=1
V1 clk avss1p8 PULSE({vdd} 0 0.0 1p 1p {Tclk/2} {Tclk}) DC 0 AC 0
V2 clr avss1p8 PULSE(0 {vdd} {-Tclk/2} 1p 1p {Tclk*2} {Tclk*30}) DC 0 AC 0
*  x1 -  4BitCounter  IS MISSING !!!!
*  x3 -  inverter  IS MISSING !!!!
C2 net2 avss1p8 1p m=1
*  x4 -  inverter  IS MISSING !!!!
C3 net3 avss1p8 1p m=1
*  x5 -  inverter  IS MISSING !!!!
C4 net4 avss1p8 1p m=1
**** begin user architecture code


* Circuit Parameters
.param vdd = 1.8
.param vss = 0.0
.param Tclk = 15n
.options TEMP = 65.0

* Include Models
.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice TT

* OP Parameters & Singals to save
.save all

* Simulations
.control
  tran 0.01u 1u
  setplot tran1
  plot clr ce+2 v(q0)+4 v(q1)+6 v(q2)+8 v(q3)+10 clk+12
reset
.endc

.end


**** end user architecture code
**.ends
.GLOBAL GND
.end
